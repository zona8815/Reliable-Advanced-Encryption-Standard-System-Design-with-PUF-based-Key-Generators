`timescale 1ns / 1ps

module Decoder(
    input [0:3] In,
    output reg [0:15] Out
);

    always@(*)begin
    
        case(In)

            4'd0 : Out = 16'b1000_0000_0000_0000;
            4'd1 : Out = 16'b0100_0000_0000_0000;
            4'd2 : Out = 16'b0010_0000_0000_0000;
            4'd3 : Out = 16'b0001_0000_0000_0000;
            4'd4 : Out = 16'b0000_1000_0000_0000;
            4'd5 : Out = 16'b0000_0100_0000_0000;
            4'd6 : Out = 16'b0000_0010_0000_0000;
            4'd7 : Out = 16'b0000_0001_0000_0000;
            4'd8 : Out = 16'b0000_0000_1000_0000;
            4'd9 : Out = 16'b0000_0000_0100_0000;
            4'd10: Out = 16'b0000_0000_0010_0000;
            4'd11: Out = 16'b0000_0000_0001_0000;
            4'd12: Out = 16'b0000_0000_0000_1000;
            4'd13: Out = 16'b0000_0000_0000_0100;
            4'd14: Out = 16'b0000_0000_0000_0010;
            4'd15: Out = 16'b0000_0000_0000_0001;
            default: Out = 16'd0;

        endcase
    
    end

endmodule